/* Custom verilog based on the template automatically generated from
/* https://wokwi.com/projects/341164910646919762 */

`ifdef SIM
`define UNIT_DELAY #1
`define FUNCTIONAL
`define USE_POWER_PINS
`include "libs.ref/sky130_fd_sc_hd/verilog/primitives.v"
`include "libs.ref/sky130_fd_sc_hd/verilog/sky130_fd_sc_hd.v"
`endif

`default_nettype none

module user_module_341164910646919762
  (
   input wire [7:0]  io_in,
   output wire [7:0] io_out
   );
   wire              clk = io_in[0];
   wire              clk_scan = io_in[1];
   wire              rstn = io_in[2];
   wire              scan_en = io_in[3];

   localparam        DIGITS = 4;
   localparam        WIDTH = 4 * DIGITS;

   wire [WIDTH-1:0]       fibonacci;

   fibonacci_341164910646919762 #(.WIDTH(WIDTH)) fib
     (.clk(clk), .rstn(rstn),
      .value(fibonacci));

   wire [3:0]             digit;

   digit_scan_341164910646919762 #(.DIGITS(DIGITS)) digit_scan
     (.clk(clk_scan), .scan_en(scan_en), .in(fibonacci),
      .out(digit));

   assign io_out[3:0] = digit;
endmodule // user_module_341164910646919762

module fibonacci_341164910646919762
  #(
    parameter WIDTH = 16
    )
   (
    input wire         clk,
    input wire         rstn,
    output wire [WIDTH-1:0] value
    );

   reg [15:0]    a;
   assign value = a;
   reg [15:0]    b;

   wire [15:0]   sum;
   adder_341164910646919762 #(.WIDTH(16)) adder
     (.a(a), .b(b), .sum(sum));

   always @(posedge clk or negedge rstn) begin
      a <= b;
      b <= sum;

      if (!rstn) begin
         a <= 1'b0;
         b <= 1'b1;
      end
   end
endmodule // fibonacci_341164910646919762

module adder_341164910646919762
  #(
    parameter WIDTH = 16
    )
   (
    input wire [WIDTH-1:0] a,
    input wire [WIDTH-1:0] b,
    output wire [WIDTH-1:0] sum
    );

   wire [WIDTH-1:0]         cout;

   sky130_fd_sc_hd__ha_1 add_first
     (.A(a[0]), .B(b[0]), .COUT(cout[0]), .SUM(sum[0]),
      .VPWR(1'b1), .VGND(1'b0));

   genvar                   i;
   generate for (i = 1; i < WIDTH; i = i + 1) begin
      sky130_fd_sc_hd__fa_1 add_rest
                     (.A(a[i]), .B(b[i]), .CIN(cout[i-1]),
                      .COUT(cout[i]), .SUM(sum[i]),
                      .VPWR(1'b1), .VGND(1'b0));
   end
   endgenerate
endmodule // adder_341164910646919762

module digit_scan_341164910646919762
  #(
    parameter DIGITS = 4
    )
   (
    input wire                clk,
    input wire                scan_en,
    input wire [4*DIGITS-1:0] in,
    output wire [3:0]         out
    );

   wire [4*DIGITS-1:0]        q;
   assign out = q[3:0];
   wire [4*DIGITS-1:0]        scd;
   assign scd = {4'b0, q[4*DIGITS-1:4]};

   genvar                     i;
   generate for (i = 0; i < 4 * DIGITS; i = i + 1) begin
      sky130_fd_sc_hd__sdfxtp_1 scan_ff
                     (.D(in[i]), .SCD(scd[i]), .SCE(scan_en),
                      .CLK(clk), .Q(q[i]),
                      .VPWR(1'b1), .VGND(1'b0));
   end
   endgenerate
endmodule // digit_scan_341164910646919762
